magic
tech scmos
timestamp 1623093546
<< nwell >>
rect -13 18 13 46
<< ntransistor >>
rect -1 7 1 12
<< ptransistor >>
rect -1 25 1 35
<< ndiffusion >>
rect -7 7 -6 12
rect -2 7 -1 12
rect 1 7 2 12
rect 6 7 7 12
<< pdiffusion >>
rect -7 25 -6 35
rect -2 25 -1 35
rect 1 25 2 35
rect 6 25 7 35
<< ndcontact >>
rect -6 7 -2 12
rect 2 7 6 12
<< pdcontact >>
rect -6 25 -2 35
rect 2 25 6 35
<< psubstratepcontact >>
rect -6 -2 -2 2
rect 2 -2 6 2
<< nsubstratencontact >>
rect -6 39 -2 43
rect 2 39 6 43
<< polysilicon >>
rect -1 35 1 37
rect -1 12 1 25
rect -1 5 1 7
<< polycontact >>
rect -5 16 -1 20
<< metal1 >>
rect -9 43 9 44
rect -9 39 -6 43
rect -2 39 2 43
rect 6 39 9 43
rect -9 38 9 39
rect -6 35 -2 38
rect -7 16 -5 20
rect 2 12 6 25
rect -6 3 -2 7
rect -9 2 9 3
rect -9 -2 -6 2
rect -2 -2 2 2
rect 6 -2 9 2
rect -9 -3 9 -2
<< labels >>
rlabel metal1 0 0 0 0 1 gnd
rlabel metal1 -6 18 -6 18 1 in
rlabel metal1 4 18 4 18 1 out
rlabel metal1 0 41 0 41 5 vdd
<< end >>
